module dcp_top();
  
endmodule
